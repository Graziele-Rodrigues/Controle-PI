library verilog;
use verilog.vl_types.all;
entity pid_vlg_vec_tst is
end pid_vlg_vec_tst;
