LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE ieee.std_logic_unsigned.all;
 
ENTITY pid IS
    PORT (
        clk: IN  STD_LOGIC; -- na placa usar 50MHz
		  enable: IN  STD_LOGIC;
		  clear: IN  STD_LOGIC;
        entrada_std : IN STD_LOGIC_VECTOR(7 DOWNTO 0); -- valor de entrada
        saida: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)  -- valor de saida
    );
	 attribute chip_pin: string;
	 attribute chip_pin of clk: signal is "N2";
	 attribute chip_pin of clear: signal is "N25";
	 attribute chip_pin of enable: signal is "N26";
	 attribute chip_pin of entrada_std: signal is "P25, AE14, AF14, AD13, AC13, B13, A13, N1";
	 attribute chip_pin of saida: signal is "AB21, AC22, AD22, AD23, AD21, AC21, AA14, Y13";
END pid;
 
ARCHITECTURE RTL OF pid IS
 
    -- valores constantes kp, ki
    constant con_kp: integer := 1;   -- Kp = 0.1 multiplicado por 10 para evitar fracoes
    constant con_kp_denominador: integer := 10;  -- Denominador para Kp
    constant con_ki: integer := 5;   -- Ki = 0.5 multiplicado por 10
    constant con_ki_denominador: integer := 10;  -- Denominador para Ki
    constant tempo_divi: integer := 1;   -- Divisor de tempo (ajustar depois)


    -- sinais internos
    signal erro_atual        : integer;
    signal erro_soma         : integer;
    signal p, i              : integer;
    signal realimentacao_reg : integer := 0;
    signal erro_soma_reg     : integer := 0;
	 signal ianterior        : integer;
	 signal integral        : integer;

 
    -- entrada / saida convertido para inteiro
    signal entrada : integer;
    signal output_val_int : integer;
	 signal output_loaded : integer;
	 
BEGIN
    -- converte entrada / saida
    entrada <= to_integer(unsigned(entrada_std));
    saida   <= std_logic_vector(to_unsigned(output_val_int, saida'length));
 
    -- calcula erros
    erro_atual       <= entrada - realimentacao_reg;
    erro_soma        <= erro_atual + erro_soma_reg;
	 
    -- calcula p 
    p <= (con_kp * erro_atual) / con_kp_denominador;
	 integral <= ianterior + erro_atual*(tempo_divi);
    -- calcula i, a parte integral, usando metodo Euler
    i <= (con_ki * integral) / con_ki_denominador;
 
    -- aplica pi
    output_loaded <= (p + i);
	
	
    PROCESS (clk)
    BEGIN
		  IF clear = '1'  THEN
				realimentacao_reg <= 0;
            output_val_int    <= 0;
            erro_soma_reg     <= 0;
				ianterior <= 0;
        ELSIF clk'event and clk = '1' and enable = '1'  THEN
				realimentacao_reg <= output_loaded;
            output_val_int    <= output_loaded;
            erro_soma_reg     <= erro_soma;
				ianterior <= integral;
        END IF;
    END PROCESS;
END RTL;